.include ibm_90nm.txt

.subckt inv 1 3 2 0
c1 3 0 10pf
MN 3 1 0 0 cmosn l=90n w=180n
MN1 3 1 2 2 cmosp l=90n w=180n
.ends

vdd 2 0 2
xinv1 4 5 2 0 inv
xinv2 5 6 2 0 inv
xinv3 6 4 2 0 inv

.control
run
tran 1n 10u
plot v(6)
.endc
.end
