.include ibm_90nm.txt

vdd 2 0 0.9
vgs 1 0 0.9
MN 2 1 0 0 cmosn l=90n w=180n

.control
run
dc vgs 0 0.9 0.01
plot log(-i(Vdd))
.endc
.end
