.include ibm_90nm.txt

c1 5 0 1pf
c2 4 0 1pf
vdd 2 0 0.9
v1 6 0 0.9

mn1 3 1 2 2 cmosp l=90n w=90n  //qbar
mn2 3 1 0 0 cmosn l=90n w=360n

mn3 1 3 2 2 cmosp l=90n w=90n  //q
mn4 1 3 0 0 cmosn l=90n w=90n

mn5 5 6 1 0 cmosn l=90n w=300n //bit
mn6 4 6 3 0 cmosn l=90n w=180n //bit bar

.ic v(5)=0.9 v(4)=0.9 v(1)=0 v(3)=0.9


.control
run
tran 1n 5u
plot v(1) v(3) v(4) v(5) 
.endc
.end
**for w/l of mn5 >320 condition fail for read
** cell ratio must be > 0.28 