.include ibm_90nm.txt

vdd 0 2 0.9
vgs 1 2 0.9
MN 0 1 2 2 cmosp l=90n w=180n

.control
run
dc vgs 0 0.9 0.01
plot log(-i(Vdd))
.endc
.end
